module features_extractor (
    
);
    
endmodule