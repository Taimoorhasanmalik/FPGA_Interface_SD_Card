module accumulator (input wire clk, reset ,input wire [7:0] data_in, input wire en, output wire [7:0] data_out);
    reg [7:0] bram [0:200];
    always @(posedge clk, posedge reset) begin
        
        
    end
    
endmodule